
/******************************************************************************
 * DVT CODE TEMPLATE: package
 * Created by serdud on Nov 2, 2023
 * amiq = amiq, ral_adapter_handshake = ral_adapter_handshake
 *******************************************************************************/

package amiq_ral_sandbox_tc_pkg;

	// UVM macros
	`include "uvm_macros.svh"
	// UVM class library compiled in a package
	import uvm_pkg::*;
	
	import amiq_ral_sandbox_env_pkg::*;
	
	`include "amiq_ral_sandbox_tc.svh"

endpackage : amiq_ral_sandbox_tc_pkg