/******************************************************************************
 * DVT CODE TEMPLATE: package
 * Created by serdud on Nov 2, 2023
 * uvc_company = amiq, uvc_name = ral_req_rsp_handshake
 *******************************************************************************/

package amiq_ral_req_rsp_handshake_pkg;

	// UVM macros
	`include "uvm_macros.svh"
	// UVM class library compiled in a package
	import uvm_pkg::*;
	
	`include "amiq_ral_req_rsp_handshake.svh"
	
endpackage : amiq_ral_req_rsp_handshake_pkg